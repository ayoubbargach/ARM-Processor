library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.instruction_field.all;

entity fetch is
  
  port (
    clk     : in std_logic;
    reset   : in std_logic;
    enable  : in std_logic;
    pc_data : in std_logic_vector(31 downto 0);
    pc_wr   : in std_logic;
    instruct_addr : out  std_logic_vector(31 downto 0);
    fetch_ok : out std_logic);

end fetch;

architecture behavioral of fetch is

  signal current_pc : unsigned(31 downto 0);
  signal pc : unsigned(31 downto 0);

begin  -- behavioral

  process(clk, reset)
  begin
    if reset = '1' then -- reset asynchrone sur niveau haut
      current_pc <= (others => '0');
      fetch_ok <= '0';
    elsif clk'event and clk = '1' then
      current_pc <= pc;
      fetch_ok <= enable;
    end if;
  end process;

  process(current_pc, pc_wr, enable)
  begin
    if pc_wr = '1' then
      instruct_addr <= pc_data;
      pc <= unsigned(pc_data);
    else
      instruct_addr <= std_logic_vector(current_pc);
      if enable = '1' then
        pc <= current_pc + 4;
      else
        pc <= current_pc;
      end if;
    end if;
  end process;

end behavioral;
